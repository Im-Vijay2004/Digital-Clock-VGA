module TITLE(clk_25MHz,title_adrs,title,name_adrs,name);
input clk_25MHz;
input [5:0] title_adrs,name_adrs;
output reg [0:499] title;
output reg [0:199] name;
always @(posedge clk_25MHz)
begin
    case(title_adrs)
        6'd00:title<=500'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd01:title<=500'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd02:title<=500'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000;
        6'd03:title<=500'b01111111111111111111110000000000000000000000000000011111110000000000000000000000000000111111111111111111000000000000000000001111111000000001111111111111111111111111111111111111100000000000000000000011111111100000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000111111111111111000000000000000001111111000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000001111111111111110000000000000000011111110000000000000000000111111100;
        6'd04:title<=500'b11111111111111111111111111000000000000000000000000011111110000000000000000000000000111111111111111111111110000000000000000001111111000000001111111111111111111111111111111111111110000000000000000000011111111100000000000000000000000000111111100000000000000000000000000000000000000000000000000000000011111111111111111111000000000000001111111000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000111111111111111111110000000000000011111110000000000000000001111111100;
        6'd05:title<=500'b11111111111111111111111111110000000000000000000000011111110000000000000000000000011111111111111111111111111100000000000000001111111000000001111111111111111111111111111111111111110000000000000000000111111111110000000000000000000000000111111100000000000000000000000000000000000000000000000000000001111111111111111111111110000000000001111111000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000011111111111111111111111100000000000011111110000000000000000011111111000;
        6'd06:title<=500'b11111111111111111111111111111100000000000000000000011111110000000000000000000000111111111111111111111111111111000000000000001111111000000001111111111111111111111111111111111111110000000000000000000111111111110000000000000000000000000111111100000000000000000000000000000000000000000000000000000111111111111111111111111111000000000001111111000000000000000000000000000000000011111111111111111111111111111100000000000000000000000001111111111111111111111111110000000000011111110000000000000000111111111000;
        6'd07:title<=500'b11111111111111111111111111111110000000000000000000011111110000000000000000000011111111111111111111111111111111100000000000001111111000000001111111111111111111111111111111111111110000000000000000001111111111110000000000000000000000000111111100000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111000000000000000000000000000000000111111111111111111111111111111110000000000000000000000011111111111111111111111111111000000000011111110000000000000000111111110000;
        6'd08:title<=500'b11111111111111111111111111111111000000000000000000011111110000000000000000000111111111111110000000011111111111100000000000001111111000000000111111111111111111111111111111111111100000000000000000001111111111111000000000000000000000000111111100000000000000000000000000000000000000000000000000011111111111111000011111111111110000000001111111000000000000000000000000000000001111111111110000000001111111111111000000000000000000000111111111111110000111111111111000000000011111110000000000000001111111100000;
        6'd09:title<=500'b11111110000000000000011111111111110000000000000000011111110000000000000000001111111111100000000000000001111111100000000000001111111000000000000000000000000111111100000000000000000000000000000000001111111111111000000000000000000000000111111100000000000000000000000000000000000000000000000000111111111110000000000001111111110000000001111111000000000000000000000000000000011111111111000000000000001111111111100000000000000000001111111111100000000000011111111100000000011111110000000000000011111111000000;
        6'd10:title<=500'b11111110000000000000000011111111110000000000000000011111110000000000000000011111111110000000000000000000011111100000000000001111111000000000000000000000000111111100000000000000000000000000000000011111111111111000000000000000000000000111111100000000000000000000000000000000000000000000000000111111111000000000000000001111110000000001111111000000000000000000000000000000111111111100000000000000000111111111100000000000000000011111111110000000000000000111111100000000011111110000000000000111111110000000;
        6'd11:title<=500'b11111110000000000000000001111111111000000000000000011111110000000000000000111111111100000000000000000000000111100000000000001111111000000000000000000000000111111100000000000000000000000000000000011111100111111100000000000000000000000111111100000000000000000000000000000000000000000000000001111111110000000000000000000111110000000001111111000000000000000000000000000000111111110000000000000000000001111111110000000000000000011111111100000000000000000001111000000000011111110000000000001111111110000000;
        6'd12:title<=500'b11111110000000000000000000011111111100000000000000011111110000000000000000111111110000000000000000000000000001100000000000001111111000000000000000000000000111111100000000000000000000000000000000011111100111111100000000000000000000000111111100000000000000000000000000000000000000000000000011111111100000000000000000000001100000000001111111000000000000000000000000000001111111100000000000000000000000111111111000000000000000111111111000000000000000000000011000000000011111110000000000001111111100000000;
        6'd13:title<=500'b11111110000000000000000000001111111110000000000000011111110000000000000001111111100000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000000111111100111111100000000000000000000000111111100000000000000000000000000000000000000000000000011111111000000000000000000000000000000000001111111000000000000000000000000000011111111100000000000000000000000011111111000000000000000111111110000000000000000000000000000000000011111110000000000011111111000000000;
        6'd14:title<=500'b11111110000000000000000000000111111110000000000000011111110000000000000011111111100000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000000111111000011111110000000000000000000000111111100000000000000000000000000000000000000000000000111111110000000000000000000000000000000000001111111000000000000000000000000000011111111000000000000000000000000011111111000000000000001111111100000000000000000000000000000000000011111110000000000111111110000000000;
        6'd15:title<=500'b11111110000000000000000000000111111111000000000000011111110000000000000011111111000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000000111111000011111110000000000000000000000111111100000000000000000000000000000000000000000000000111111110000000000000000000000000000000000001111111000000000000000000000000000011111110000000000000000000000000001111111100000000000001111111000000000000000000000000000000000000011111110000000001111111100000000000;
        6'd16:title<=500'b11111110000000000000000000000011111111000000000000011111110000000000000111111110000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000001111111000011111111000000000000000000000111111100000000000000000000000000000000000000000000001111111100000000000000000000000000000000000001111111000000000000000000000000000111111110000000000000000000000000001111111100000000000011111111000000000000000000000000000000000000011111110000000011111111000000000000;
        6'd17:title<=500'b11111110000000000000000000000001111111100000000000011111110000000000000111111110000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000001111110000001111111000000000000000000000111111100000000000000000000000000000000000000000000001111111000000000000000000000000000000000000001111111000000000000000000000000000111111100000000000000000000000000000111111110000000000011111110000000000000000000000000000000000000011111110000000011111111000000000000;
        6'd18:title<=500'b11111110000000000000000000000001111111100000000000011111110000000000001111111100000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000001111110000001111111000000000000000000000111111100000000000000000000000000000000000000000000011111111000000000000000000000000000000000000001111111000000000000000000000000001111111100000000000000000000000000000111111110000000000111111110000000000000000000000000000000000000011111110000000111111110000000000000;
        6'd19:title<=500'b11111110000000000000000000000001111111100000000000011111110000000000001111111100000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000011111110000001111111100000000000000000000111111100000000000000000000000000000000000000000000011111111000000000000000000000000000000000000001111111000000000000000000000000001111111100000000000000000000000000000111111110000000000111111110000000000000000000000000000000000000011111110000001111111100000000000000;
        6'd20:title<=500'b11111110000000000000000000000000111111100000000000011111110000000000001111111000000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000011111100000000111111100000000000000000000111111100000000000000000000000000000000000000000000011111110000000000000000000000000000000000000001111111000000000000000000000000001111111000000000000000000000000000000011111110000000000111111100000000000000000000000000000000000000011111110000011111111000000000000000;
        6'd21:title<=500'b11111110000000000000000000000000111111110000000000011111110000000000011111111000000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000111111100000000111111100000000000000000000111111100000000000000000000000000000000000000000000011111110000000000000000000000000000000000000001111111000000000000000000000000001111111000000000000000000000000000000011111110000000000111111100000000000000000000000000000000000000011111110000111111110000000000000000;
        6'd22:title<=500'b11111110000000000000000000000000111111110000000000011111110000000000011111111000000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000111111100000000111111110000000000000000000111111100000000000000000000000000000000000000000000011111110000000000000000000000000000000000000001111111000000000000000000000000001111111000000000000000000000000000000011111110000000001111111100000000000000000000000000000000000000011111110000111111100000000000000000;
        6'd23:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111111000000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000000111111000000000011111110000000000000000000111111100000000000000000000000000000000000000000000111111110000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000000000000011111111000000001111111100000000000000000000000000000000000000011111110001111111100000000000000000;
        6'd24:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111110000000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000001111111000000000011111110000000000000000000111111100000000000000000000000000000000000000000000111111110000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000000000000011111111000000001111111100000000000000000000000000000000000000011111110011111111000000000000000000;
        6'd25:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111110000000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000001111111000000000001111111000000000000000000111111100000000000000000000000000000000000000000000111111110000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000000000000011111111000000001111111000000000000000000000000000000000000000011111110111111110000000000000000000;
        6'd26:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111110000000000000000000000000000000000000000000000001111111000000000000000000000000111111100000000000000000000000000001111110000000000001111111000000000000000000111111100000000000000000000000000000000000000000000111111100000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000000000000011111111000000001111111000000000000000000000000000000000000000011111111111111100000000000000000000;
        6'd27:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111110000000000000001111111111111111111000000000000001111111000000000000000000000000111111100000000000000000000000000011111110000000000001111111100000000000000000111111100000000000000000000000000000000000000000000111111100000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000000000000011111111000000001111111000000000000000000000000000000000000000011111111111111100000000000000000000;
        6'd28:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111110000000000000001111111111111111111100000000000001111111000000000000000000000000111111100000000000000000000000000011111110000000000000111111100000000000000000111111100000000000000000000000000000000000000000000111111100000000000000000000000000000000000000001111111000000000000000000000000011111110000000000000000000000000000000011111111000000001111111000000000000000000000000000000000000000011111111111111110000000000000000000;
        6'd29:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111110000000000000001111111111111111111100000000000001111111000000000000000000000000111111100000000000000000000000000011111100000000000000111111100000000000000000111111100000000000000000000000000000000000000000000111111100000000000000000000000000000000000000001111111000000000000000000000000011111110000000000000000000000000000000011111111000000001111111000000000000000000000000000000000000000011111110111111110000000000000000000;
        6'd30:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111110000000000000001111111111111111111100000000000001111111000000000000000000000000111111100000000000000000000000000111111100000000000000111111110000000000000000111111100000000000000000000000000000000000000000000111111100000000000000000000000000000000000000001111111000000000000000000000000011111110000000000000000000000000000000011111111000000001111111000000000000000000000000000000000000000011111110011111111000000000000000000;
        6'd31:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111110000000000000001111111111111111111100000000000001111111000000000000000000000000111111100000000000000000000000000111111100000000000000011111110000000000000000111111100000000000000000000000000000000000000000000111111100000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000000000000011111111000000001111111000000000000000000000000000000000000000011111110011111111100000000000000000;
        6'd32:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111110000000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000000001111111000000000000000011111110000000000000000111111100000000000000000000000000000000000000000000111111110000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000000000000011111111000000001111111000000000000000000000000000000000000000011111110001111111110000000000000000;
        6'd33:title<=500'b11111110000000000000000000000000011111110000000000011111110000000000011111110000000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000000001111111000000000000000011111111000000000000000111111100000000000000000000000000000000000000000000111111110000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000000000000011111111000000001111111000000000000000000000000000000000000000011111110000111111110000000000000000;
        6'd34:title<=500'b11111110000000000000000000000000111111110000000000011111110000000000011111110000000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000000001111110000000000000000001111111000000000000000111111100000000000000000000000000000000000000000000111111110000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000000000000011111110000000001111111100000000000000000000000000000000000000011111110000011111111000000000000000;
        6'd35:title<=500'b11111110000000000000000000000000111111110000000000011111110000000000011111111000000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000000011111111000000000000000001111111000000000000000111111100000000000000000000000000000000000000000000111111110000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000000000000011111110000000001111111100000000000000000000000000000000000000011111110000011111111100000000000000;
        6'd36:title<=500'b11111110000000000000000000000000111111110000000000011111110000000000011111111000000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000000011111111111111111111111111111111100000000000000111111100000000000000000000000000000000000000000000011111110000000000000000000000000000000000000001111111000000000000000000000000001111111000000000000000000000000000000011111110000000001111111100000000000000000000000000000000000000011111110000001111111110000000000000;
        6'd37:title<=500'b11111110000000000000000000000000111111100000000000011111110000000000011111111000000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000000011111111111111111111111111111111100000000000000111111100000000000000000000000000000000000000000000011111110000000000000000000000000000000000000001111111000000000000000000000000001111111000000000000000000000000000000011111110000000000111111100000000000000000000000000000000000000011111110000000111111110000000000000;
        6'd38:title<=500'b11111110000000000000000000000001111111100000000000011111110000000000001111111100000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000000111111111111111111111111111111111100000000000000111111100000000000000000000000000000000000000000000011111111000000000000000000000000000000000000001111111000000000000000000000000001111111100000000000000000000000000000111111110000000000111111100000000000000000000000000000000000000011111110000000011111111000000000000;
        6'd39:title<=500'b11111110000000000000000000000001111111100000000000011111110000000000001111111100000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000000111111111111111111111111111111111110000000000000111111100000000000000000000000000000000000000000000011111111000000000000000000000000000000000000001111111000000000000000000000000001111111100000000000000000000000000000111111100000000000111111110000000000000000000000000000000000000011111110000000011111111100000000000;
        6'd40:title<=500'b11111110000000000000000000000001111111000000000000011111110000000000001111111110000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000000111111111111111111111111111111111110000000000000111111100000000000000000000000000000000000000000000011111111000000000000000000000000000000000000001111111000000000000000000000000001111111100000000000000000000000000000111111100000000000111111110000000000000000000000000000000000000011111110000000001111111110000000000;
        6'd41:title<=500'b11111110000000000000000000000011111111000000000000011111110000000000000111111110000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000001111111100000000000000000000111111111000000000000111111100000000000000000000000000000000000000000000001111111100000000000000000000000000000000000001111111000000000000000000000000000111111110000000000000000000000000001111111100000000000011111111000000000000000000000000000000000000011111110000000000111111110000000000;
        6'd42:title<=500'b11111110000000000000000000000011111111000000000000011111110000000000000111111111000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000001111111000000000000000000000011111111000000000000111111100000000000000000000000000000000000000000000001111111100000000000000000000000000000000000001111111000000000000000000000000000111111110000000000000000000000000001111111000000000000011111111000000000000000000000000000000000000011111110000000000011111111000000000;
        6'd43:title<=500'b11111110000000000000000000000111111110000000000000011111110000000000000011111111000000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000011111111000000000000000000000001111111000000000000111111100000000000000000000000000000000000000000000000111111110000000000000000000000000000000000001111111000000000000000000000000000111111111000000000000000000000000011111111000000000000011111111100000000000000000000000000000000000011111110000000000011111111100000000;
        6'd44:title<=500'b11111110000000000000000000001111111110000000000000011111110000000000000011111111100000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000011111110000000000000000000000001111111100000000000111111100000000000000000000000000000000000000000000000111111111000000000000000000000000000000000001111111000000000000000000000000000011111111000000000000000000000000111111110000000000000001111111100000000000000000000000000000000000011111110000000000001111111110000000;
        6'd45:title<=500'b11111110000000000000000000011111111100000000000000011111110000000000000001111111110000000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000011111110000000000000000000000001111111100000000000111111100000000000000000000000000000000000000000000000111111111000000000000000000000001110000000001111111000000000000000000000000000011111111100000000000000000000001111111110000000000000001111111110000000000000000000000011100000000011111110000000000000111111110000000;
        6'd46:title<=500'b11111110000000000000000000111111111000000000000000011111110000000000000000111111111100000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000111111110000000000000000000000000111111100000000000111111100000000000000000000000000000000000000000000000011111111110000000000000000000011110000000001111111000000000000000000000000000001111111110000000000000000000011111111100000000000000000111111111000000000000000000001111100000000011111110000000000000011111111000000;
        6'd47:title<=500'b11111110000000000000000011111111110000000000000000011111110000000000000000011111111110000000000000000000111111100000000000001111111000000000000000000000000111111100000000000000000000111111100000000000000000000000000111111110000000000111111100000000000000000000000000000000000000000000000001111111111000000000000000001111110000000001111111000000000000000000000000000000111111111000000000000000000111111111100000000000000000011111111110000000000000000011111100000000011111110000000000000011111111100000;
        6'd48:title<=500'b11111110000000000000011111111111100000000000000000011111110000000000000000011111111111100000000000000011111111100000000000001111111000000000000000000000000111111100000000000000000000111111100000000000000000000000000111111110000000000111111110000000000000000000000000000000000000000000000000111111111110000000000001111111110000000001111111000000000000000000000000000000111111111110000000000000011111111111000000000000000000011111111111100000000000011111111100000000011111110000000000000001111111110000;
        6'd49:title<=500'b11111111111111111111111111111111000000000000000000011111110000000000000000001111111111111111000000111111111111100000000000001111111000000000000000000000000111111100000000000000000001111111000000000000000000000000000011111110000000000111111111111111111111111111000000000000000000000000000000111111111111111100011111111111110000000001111111111111111111111111110000000000011111111111110000000011111111111110000000000000000000001111111111111111000111111111111100000000011111110000000000000000111111110000;
        6'd50:title<=500'b11111111111111111111111111111110000000000000000000011111110000000000000000000011111111111111111111111111111111100000000000001111111000000000000000000000000111111100000000000000000001111111000000000000000000000000000011111111000000000111111111111111111111111111000000000000000000000000000000011111111111111111111111111111100000000001111111111111111111111111110000000000001111111111111111111111111111111100000000000000000000000111111111111111111111111111111000000000011111110000000000000000011111111000;
        6'd51:title<=500'b11111111111111111111111111111100000000000000000000011111110000000000000000000001111111111111111111111111111111000000000000001111111000000000000000000000000111111100000000000000000001111111000000000000000000000000000001111111000000000111111111111111111111111111000000000000000000000000000000000111111111111111111111111111000000000001111111111111111111111111110000000000000111111111111111111111111111111000000000000000000000000011111111111111111111111111110000000000011111110000000000000000011111111100;
        6'd52:title<=500'b11111111111111111111111111110000000000000000000000011111110000000000000000000000011111111111111111111111111110000000000000001111111000000000000000000000000111111100000000000000000011111110000000000000000000000000000001111111100000000111111111111111111111111111100000000000000000000000000000000011111111111111111111111110000000000001111111111111111111111111110000000000000001111111111111111111111111100000000000000000000000000000111111111111111111111111100000000000011111110000000000000000001111111100;
        6'd53:title<=500'b11111111111111111111111110000000000000000000000000011111110000000000000000000000000111111111111111111111111000000000000000001111111000000000000000000000000111111100000000000000000011111110000000000000000000000000000001111111100000000011111111111111111111111111000000000000000000000000000000000000111111111111111111111000000000000001111111111111111111111111110000000000000000011111111111111111111110000000000000000000000000000000001111111111111111111110000000000000011111110000000000000000000111111110;
        6'd54:title<=500'b01111111111111111111100000000000000000000000000000011111110000000000000000000000000001111111111111111111000000000000000000001111111000000000000000000000000111111100000000000000000011111110000000000000000000000000000000111111100000000011111111111111111111111111000000000000000000000000000000000000001111111111111111000000000000000000111111111111111111111111110000000000000000000111111111111111111000000000000000000000000000000000000011111111111111110000000000000000011111110000000000000000000011111110;
        6'd55:title<=500'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000;
        6'd56:title<=500'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6'd57:title<=500'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        default:
                title<=500'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
end
always @(posedge clk_25MHz)
begin
    case(name_adrs)
    6'd00:name<=200'b00111000000000001110000000001111111111110000000110000000001110011000000011000000001110000000110000000110000000111000000001110000000010000011111111000000001100000000110000111111110000000000111000000000;
    6'd01:name<=200'b00111100000000001110000000001111111111110000000110000000001100011000000011000000001110000000110000001110000001111000000001111000000110000011111111110000001100000000110000111111111000000000111100000000;
    6'd02:name<=200'b00111100000000011110000000000000011000000000000111000000001100011000000011000000011111000000111000001100000001111000000001111100000110000011000000111000001100000000110000110000011100000000111100000000;
    6'd03:name<=200'b00111110000000011110000000000000011000000000000011000000011100011000000011000000011011000000011000011100000001101100000001101100000110000011000000011100001100000000110000110000001100000001101100000000;
    6'd04:name<=200'b00110110000000110110000000000000011000000000000011000000011000011000000011000000011011000000011100011000000011001100000001101110000110000011000000001100001100000000110000110000001100000001101110000000;
    6'd05:name<=200'b00110110000000110110000000000000011000000000000011100000011000011000000011000000110001100000001100011000000011001110000001100110000110000011000000001100001100000000110000110000001100000011000110000000;
    6'd06:name<=200'b00110011000001100110000000000000011000000000000001100000110000011000000011000000110001100000001110111000000011000110000001100111000110000011000000001100001100000000110000110000011100000011000110000000;
    6'd07:name<=200'b00110011000001100110000000000000011000000000000001100000110000011000000011000001110001110000000111110000000110000110000001100011000110000011000000001110001111111111110000111111111000000011000111000000;
    6'd08:name<=200'b00110011100001100110000000000000011000000000000000110000110000011000000011000001100000110000000011110000000110000111000001100011100110000011000000001110001111111111110000111111110000000110000011000000;
    6'd09:name<=200'b00110001100011000110000000000000011000000000000000110001100000011000000011000001100000110000000011110000000110000011000001100001100110000011000000001110001100000000110000110001110000000110000011000000;
    6'd10:name<=200'b00110001100011000110000000000000011000000000000000110001100000011000000011000011111111111000000001100000001111111111000001100000110110000011000000001100001100000000110000110000011000000111111111100000;
    6'd11:name<=200'b00110000110110000110000000000000011000000000000000011001100000011000000011000011111111111000000001100000001111111111100001100000110110000011000000001100001100000000110000110000011000001111111111100000;
    6'd12:name<=200'b00110000110110000110000000000000011000000000000000011011000000011000000011000011000000011000000001100000011100000001100001100000011110000011000000011100001100000000110000110000011100001100000001110000;
    6'd13:name<=200'b00110000111110000110000000000000011000000000000000011111000000011000000011000111000000011100000001100000011000000001100001100000011110000011000000111000001100000000110000110000001100001100000000110000;
    6'd14:name<=200'b00110000011100000110000000000000011000000000000000001111000000011000100111000110000000001100000001100000011000000001110001100000001110000011000011110000001100000000110000110000001110011000000000110000;
    6'd15:name<=200'b00110000011100000110000000000000011000000000000000001110000000011000111110000110000000001100000001100000111000000000110001100000001110000011111111100000001100000000110000110000000110011000000000111000;
    6'd16:name<=200'b00110000001000000110000000000000000000000000000000000100000000001000011100000100000000000100000001100000010000000000010000000000000010000001111000000000000000000000100000010000000000010000000000010000;
    6'd17:name<=200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    6'd18:name<=200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    6'd19:name<=200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    6'd20:name<=200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    6'd21:name<=200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    6'd22:name<=200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    6'd23:name<=200'b00000011111000000000000001100000000000011000000000111111000000001100000000100000110011111111111110011000000001100000000001100000001000011000000001100000111000000000000110000000001100000000001111100000;
    6'd24:name<=200'b00001111111110000000000011110000000000111100000011111111100000001100000001100000110011111111111110011000000001100000000001100000011000011000000001100000111100000000001110000000001110000000011111111000;
    6'd25:name<=200'b00011100000111000000000011110000000000111100000111000001110000001100000001100000110000000011000000011000000001100000000001100000111000011000000001100000111100000000011110000000011110000000011000011100;
    6'd26:name<=200'b00111000000000000000000011011000000001101100000110000000111000001100000001100000110000000011000000011000000001100000000001100001110000011000000001100000111100000000011110000000011111000000011000001110;
    6'd27:name<=200'b00110000000000000000000011011000000001101100001110000000011100001100000001100000110000000011000000011000000001100000000001100011100000011000000001100000110110000000110110000000110011000000011000000110;
    6'd28:name<=200'b01110000000000000000000011011100000011001100001100000000011100001100000001100000110000000011000000011000000001100000000001100011000000011000000001100000110110000000110110000000110011000000011000000110;
    6'd29:name<=200'b01100000000000000000000011001100000011001100001100000000001100001100000001100000110000000011000000011000000001100000000001100110000000011000000001100000110111000000110110000000110011100000011000001110;
    6'd30:name<=200'b01100000000000000000000011001100000011001100011100000000001100001111111111100000110000000011000000011111111111100000000001111100000000011000000001100000110011000001100110000001100001100000011000011100;
    6'd31:name<=200'b01100000111111000000000011000110000110001100011100000000001100001111111111100000110000000011000000011111111111100000000001111100000000011000000001100000110011000001100110000001100001100000011111111000;
    6'd32:name<=200'b01100000111111000000000011000110000110001100011100000000001100001100000001100000110000000011000000011100000001100000000001111110000000011000000001100000110001100011000110000001100000110000011111111000;
    6'd33:name<=200'b01100000000011000000000011000111001100001100011100000000001100001100000001100000110000000011000000011000000001100000000001100111000000011000000001100000110001100011000110000011000000110000011000011000;
    6'd34:name<=200'b01100000000011000000000011000011001100001100001100000000011100001100000001100000110000000011000000011000000001100000000001100011000000011000000001100000110001110111000110000011111111111000011000001100;
    6'd35:name<=200'b01110000000011000000000011000011011100001100001100000000011000001100000001100000110000000011000000011000000001100000000001100001100000011000000001100000110000110110000110000011111111111000011000001100;
    6'd36:name<=200'b00111000000011000000000011000001111000001100001110000000011000001100000001100000110000000011000000011000000001100000000001100001110000011100000011100000110000111110000110000110000000011000011000000110;
    6'd37:name<=200'b00111100000011000000000011000001111000001100000111000001110000001100000001100000110000000011000000011000000001100000000001100000111000001100000011000000110000011100000110000110000000011100011000000110;
    6'd38:name<=200'b00011111111111000000000011000001110000001100000011111111110000001100000001100000110000000011000000011000000001100000000001100000011000001111111111000000110000011100000110001110000000001100011000000110;
    6'd39:name<=200'b00000111111100000000000011000000110000001100000001111111000000001100000001100000110000000011000000011000000001100000000001100000001100000011111100000000110000011000000110001100000000001100011000000110;
    endcase
end
endmodule